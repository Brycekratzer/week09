module dLatch (
    input D, E,
    output Q,Qn
);
    @always(D,E)begin
        if()
    end
endmodule