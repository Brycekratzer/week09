module memblock8bit(
    input [7:0]InputData,
    input E,
    output [7:0]OutputData,
);

endmodule